    localparam FETCH = 8'h0;
    localparam NOP = 8'h3;
    localparam ILLEGAL = 8'h4;
    localparam UNIMP = 8'h6;
    localparam INIT_PC = 8'h7;
    localparam LW = 8'h8;
    localparam SW = 8'hd;
    localparam LB = 8'h12;
    localparam SB = 8'h17;
    localparam LH = 8'h1c;
    localparam SH = 8'h21;
    localparam LBU = 8'h26;
    localparam LHU = 8'h2b;
    localparam LUI = 8'h30;
    localparam ADDI = 8'h31;
    localparam SLTI = 8'h34;
    localparam SLTIU = 8'h37;
    localparam SLLI = 8'h3a;
    localparam SRLI = 8'h3d;
    localparam SRAI = 8'h40;
    localparam ANDI = 8'h43;
    localparam ORI = 8'h46;
    localparam XORI = 8'h49;
    localparam ADD = 8'h4c;
    localparam SUB = 8'h4f;
    localparam SLT = 8'h52;
    localparam SLTU = 8'h55;
    localparam SLL = 8'h58;
    localparam SRL = 8'h5b;
    localparam SRA = 8'h5e;
    localparam AND = 8'h61;
    localparam OR = 8'h64;
    localparam XOR = 8'h67;
    localparam JAL = 8'h6a;
    localparam JALR = 8'h6f;
    localparam AUIPC = 8'h74;
    localparam BEQ = 8'h78;
    localparam BNE = 8'h7c;
    localparam BLT = 8'h80;
    localparam BLTU = 8'h85;
    localparam BGE = 8'h8a;
    localparam BGEU = 8'h8f;
    localparam BZ_TAKEN = 8'h94;
    localparam CSRRW = 8'h98;
    localparam CSRRC = 8'h9d;
    localparam CSRRS = 8'ha2;
    localparam CSRRWI = 8'ha7;
    localparam CSRRCI = 8'hac;
    localparam CSRRSI = 8'hb1;
    localparam DRET = 8'hb6;
    localparam MRET = 8'hb6;
    localparam ECALL = 8'hb6;
    localparam EBREAK = 8'hb6;
    localparam WFI = 8'hb8;
    localparam EHALT = 8'hb9;
    localparam EXTRA = 8'hba;
